�io���\��������:8[9U6�^�$��9^���2ឡ<Q����Ϫ������ҳ&�:!qڨ���<�^@Ϭ��'�<��
��oR�4�\dl��n�W�OђD��g�A[�G�])�*����y�.!.��Y��K
Է�4��3fM��N��GG����?����� *�@��,��)���Xxg^6����s�VF�݅&cHJ��*{�U/~ݦ$}��uύ����,�}������:Á�W`>��RF��b����k�[���b
ҽ�!ՎeF�'�����|�jٻbh>��C��~P��ϛ���-����4)��v���
�ɽ'�> -(tS���Zˇ}!��w&�����.;h����)mа9��37mU,{�	��9�Qw���G�I�zX�PT�}"oo[�����`XK��÷�Tt��(\RT�v
�m��_9*��n�j��hA�.���'/�D T{O�#��4�P���`l��,Z1�"���5��7>�2��R	�����|ys畑ׁ�N�Z\O� r��p-=��U�^�+j���=��:�%U���B���u<�~ȏ����?D[�S����KȖ92A� �\�+�(W����y�J/�?ٷW���?��%�>'���k�1C">9�AY��9����R5�o�sr�+(��=�7��*�Hx�7�{�YN����:�}12*?�r�H^D��48ڸ���=L���R�>mS�)���˚�񕗘,�d���n[е����!Zh����-�@�ϔ��4�%[���Ǔ�=�� �e���̢�)��,��·�K�Ar�`�b_��0���Ϟh�`����Uɍ9|o+��B�S-+�KN	�G�j�.���@����Lp}�k�4�I��ٷ��dPY�V��x�n�'n(\I~6цIeM1t̐��(�Z�At�ء������\����x�}�ԡ,6l��H��W#�;$����٫����_HӃ��,�w�i�I�u�d��Eg�K*���¡Ah��u�2`6�[5ՙ�-th�W�T�)���{r}/[I����[cÐkѹ�:��ˊ�Ա�,�j��y�,e�L��O=��guDS2��o�h���,�SRco����b4ˢ�Ĳ��h7<��!u�6G.�ه:*	R���G���ox�k��u�<�<�3�0��p~w�?�N�$(s\uh�2y?��I���9&A>ͬ�z��<�MJ���b��<�y���[͈�� O��>�懆�zUXm��⮇�0����&1�s>ߚ>�_~8 �S�v��\}����Iڰha���x5��L�/S`�c\�|�3i��ž�N�"�W��\�Y�]0��ĩh��|-Ω���SS��]PV^HyۀoO�
��b1:��j��Z&m�������)׫�DP;䄨ȋD�pr�v�fUU��9�&;b�ra���dѹ���j7��2 1-^�k|h�o&��(���^TU�R&���=�(UY�'"/͏��Ypʿ{D�8"�aWH�f�Ӽ3_�(:���lS!R�����u!U� ۻ�����ӗ��,+���j'%�8/����4!�9[�;�!��믿~����jL�j8L��\�MLуO(֒h{�.�p�P��\�-Gћ�܈�u268E�����]>����s& ���|���hV�@�gNu��Q�x3@F�D���9��N��m���w6Ƒ��c��AoX��q�1Q�{��xBLz�u�"�
�C$�ۍ21���%�n�Ȗ�oKO&pvy�[���mJ?V��i�ǔN҇Wxa����fP�lB~�Ws�Q�9�y�HD�y�pV�B��W��̧'I��a���_}G�ҷ��+b�[���XH�$�s2��"a��� ��s�
�Q��5C^2/��r�i�[��:�I�ϊI�fKr{kmq���nMiQ3�@')��kw�&厛����4��_9:��	�Ɠ�gIQ�Ex�_a����o�b��~�JM������7�x��}�
s *��ߍ܏:����G+t�:g?�ХCt��EJv��!���<��`��.�w|�ao��}�sG�z���D�I�9균G�l�����\"�h�S���h�֞sz��"���>E��E\�E���^l�6D��̬Ȯ��_���� z�L�\�r�l��c����FC�ֶ�	_]~ف'��!�r_���g>�H����1��_%5�й(X?���
9�>����-�3�xsٗ�K�ђ�R����֏>\�4��]����cbE�y�>�^�BSBt�T�ye����\�ݗ��/]r��N�)�϶���氛� q��R���5c>l��Ј�U��Q�
��*�~�&:�uv3�y�{� �=�9��JՈ\͔���π�δ�����՟���n^Aܬ5�ތ<6˓it��5Dۆ��w����Ғᨹ/��,�Z����
])������4'�*9SҠ��w{�T.��Sz#R�j�Lܻx6�$n��R '#}�2J��fQ�ے���6s�}��}�%�#�䎮5����'�jA\;�Dp�Z��Z��F���w�/�q.u�D�̣ǰI�ZLJIv��ɧ���I5woc��:��Ԩ�n��V�МK��4o������7�p��l����G����R%���3�[Y��]��d�+�wrb�~8I�G���m�W������p���YҍwF�������L�N�x��J��p/�u.�Ê�	����A0zR!@3���)lx�	]$�@���1�K��\=����m9��0"��3�X��Ʊ��*k�uJ둑�����R�I���Qy���Z��&����0a�>�w�x�����D���ґ��J[&��x���&�	�o���Q��8�����H⬑)lx��B���Q��AU�Y�H��Y��@�Ƞ����ƣ�+�̓����IP�"zn�)���l�dG3|�*.*Zf�ճLڃ��&%����1V�O!������-���g�o��F�U�jc\V�qMEׁ���ěR� &��u��yG���v�e��l��_�2��:`��
u!>}$����X�*?�2�!�|�r�2�u����޼��9��ͫy�����>p=��[7�㉌��9��w*Z,�ƣ!�B5�O�n��J��?>�SҚ�Q�ɐ�ޭL�7LɻT�{[u/���ٻ��-��	s�����I���Jj#Fdam%�\Gt��F�C�h�Ŭ��L3�U���.�&�����~V���E��49��:<�g\1)�r�Q����Y��1m��Rڡ�5qx+�u�h��o�� 8���{�-�[EA�Оo2�{2y2�N2�K��:�1�q����RG�UQ�x�xu�9�!����g��?&�0ǝ��*�[��n}����y�q_d{_��F{Co���)]�,�5
��������J��,��c	1�2� u����a%H=��$�Db�7kډ�k�ݚh�A*�|S��4q�l�/3�kui;fN5�n|�5�S;�eB���2�_k��+��x{�s+;��:<̌��m�����P�E�R�#H��"�4G�[̑
W��n�1W��s��pМ�<�T5��/ ��s��Y�z�! f��G�|z�Oc�΃nn�!P��w�v���T&�_�)��"�(6kQ~T	��n79�a�Ԕ/���+��a�_U�jB�;����!����hc������5��{���ݟ��3eu8���$COM�:��o2|���JU���o���`np��85#��yb'겢�ݰY��X9��Vkk�ɴ�� P��[�fc��A۶�&.�����Q�]?�����|矕�o;��@����%��gAcJ�� �N��f��ꊇK�o�ȇJ+��E�]����ӥӔp�L�>E)3�T��5f�����P��*z�粐
F �>e��ݨ�6�p���~��証4:�=nN���}3q����vN;QO�e��u�Qo�w�aiUfN���	�1�� *�'���z�߮c�FH�R1[�_MZ�7TA"�%qN�T>,޷4�(*(���T,��|�1LX�I��-'���摲�>}W��� �Jш�]arx�Q1/!!�3ޝ�ŭ�I�"�Z�EuK��g]�ľ��Mj�s9�	�#�Pþ��$+<����0����rI����L��/5��ZGL�G���.ⵀr�M_���Y{H~�<��̟���L>� ��M]`tO�ۤƪ�X<�0(��E����r`�>I��p7K��6c�W�����6e�Ԑ�}A	i�ܙ	�M��*�\�s��aݐ&���1tл2��"e��p�4���x��5$��/<wkJcr1�`�#�����=X��ٕD1��CH�����qW�������/T`���\�/H�"4^=M���qܫ���o;�h��P�&S��yjiU]��m�u�]݊�.��;׏R���D��曜r��D�6A��ݎ]�Kh+�B��3��Z�cA~K��雠[1��m�v�îԗQ�M@���%(�q���W*e�~��|�->Bi�ܬM��v�����C���#_����eҥݪ���#��q�ۊ����0�zC���On��H団�=��}_���G^K\����V���2&���]cQ��k�c_��w�0�z+^��A��V�ѳ� ���i[7�����H�u����������%)�ڳ�~���:��t����{�ra���X��m\�5ȧ��,-޽�S��+�
�ԝ'	�;.7�V����zh�iw:� ��䦺�!�����}��5������ݛ�#�‌�K�x�V�m�����1�I�l��l����_��8�f\{X�""6�r|�@�%�����
N����HI�io:�<z�,�?��0Ҹ��?.�9)!�D�E��Q[��A�0��P'���0��zl�K`���tڕ-.IuhMi�U�bd�ɫ���x^.��)ɺJ�X�덬�0-��F觞�j�)��`�hg"
Ek�L��HV�fGW�^%whK��f��,�u0󚟥\T��3b�� �h&cuʟ�����:b���pNPR-���;��)2�Gm�m2�1Ǣ�ʂ[���E���T` �!�(�_��-�&"w$�hK{���R���Xx0N�t��A��P�U;&����7����v
q�8��@�Z�����[ ��6L{�9���*KA"��K������o$� ���w�5M�b�FH��E�߸ ��9��"+8���vB&T��z�9�k��y��mgCn�vm���v��ou#��0ѣ]�DkPQZV��$�C��ɻ�d@S� ]52���JvdL�"�Q�Ѐ��W�P~aG`�R�@SfUX�m�vp/be��|��=4Ӏf��هo������;o��"q��Ck���c��{�������7�'qT�����!� �����V5����'�g��|����B��@���� �WfÕ���`�/|a�v�LH��.C�ܶ���t�� 6��bI��'`p�Vŷ���3$��`�C�C�����~�	��_�O���I��!"�~��'#z��T��ɠ]L��n�c�
5�rQz�O�S�*#'�[m?�������C��@-���R`̰o����TɕB؝+4$ӆܔ��w��T R&�� {��Vm�1��H��Ԇ��>��;�P˨��\X�&�埿�[d��h��-��z7C5�������	�Ŏc
��j�DxP�@���pC�#qq]�,آ���n�a���ɓ�!#TNƤ�u�o�� ���UGa��8��&cU,׶5]OJe|���53� }S�'�<qz �o8��})wp���dK���$+���
}H��;1�����̻BŧWQ��C�:6<����D��w�@p4��i���b>�f;
K�1ױ�^���J'%/�4&�ps�e��{-�C���_D=��e�K!�id#��j%��T���Z��������O�{�iE�W���-&HC������ ��f��ڙK0�3mH�B)6՝���ۊ�I3j	�h�����8߲ϼp�uQi��&��?7	���E�c�ų\��ɜ��GDϕ�>�1=;ފC>�~Rm̯��w,�5Q��r+�c�W�Rm�p�J�M�[@�#ǐe�
���S�'lK��'��GW������*����b�#���,]�O�����.�2[��v�L���G���$!-��|���K�aڨ�'�zS���`���F���`��Mt��앫��w7���F,�s�Փ�31q76�(iHMȇ����G�6Y���A}1O�M�}�Z�.U6Y�:�w�IZ*�μ)w�zW
���mw�b[���Wʭ����t6����(��c��ɥt�b�E�37q�?���ML��*`<<DY��D�)|%�G�d]B���aC���V7$�����׀s*�q᱑�v�e��a^�U�H-�LT�6)ˡ�]s��(g��M,,�v�(���a�3�p�?i�ɸ$�6n:����xH����6��4�i�v	�A|��^~\��0�i2w���n<�Ƭ� �0�p��'њ����g�$ܢ��)m �`��@U�x9��#����k�*�^����\쩴��v��/1�� �8
��"�����b {E�%�b����ղ��B��D�͏��a?]���}�En��7��q�$ R�͑?n��Հ��1�t2rL��1��£��1λ?T*h�P�۰؎�n(*4|�e*��e�7����K=6�zK*�"��[!$@��.��>��s'ߊ��0@.'զ����<��3����)���	��A��b�Z�~{�wA0*
��mLR� ¥�M�D\�<oi���͒I�Ԅ	@@�%��'�ξ�[���1�ll�����5���a����m��JR3M�&!ր0!�5�Χ�%J��58�M�_-B3 �n2Ƙ(�#FU�ctw��H�B0�l�S����;ghw
���	�dF��?1J��$n�"�:��@�[�>��K
