"K��|�����jJ� xV;�8��~������or6'm��k�+�(30��	|;@�"�w�����ND�)�A��i��R�K��Aޚ����e`:�4��3�|t�d����q,�X.'��Զ;��8�d�'����4z�[��Bm%�4;�U���F���KW�}i=�>o��YQ��{b���vZ-yO���T=����9��FݐvZ��8K��mf��f�?���X�|�"�������^�v�ӏF��7ZA��:S]�pNν��^��h��D�k�(��bn�8���~"�bW:��=�bk��Ib���8
�:���n-֌B@cA!z~w��J�@;F^+O&QI�0�0�;�@�����J�F�2�U�/���фw�&�-꓊V#�c|~ӕQ�>}p��%�.'�D�lwf��F�rՃ��Z�;~R<vP�['����֚Xɵ���o�/�x��( ��Pl�Ɛ�;!G��@@��f\��{LV��s����@���~� K�:�&	b��ΐ��~v?�(Z}�e���1��-�~0�����rQ�� ��=�WL���������2Yԁ`L߻����[Fưz2����c��f�yU�1�.чmB�&��\���\�� ���Q)�V>W��G[��$%;�����
Q��G�ƤG,g����n�	�lY/��!7j_��À���7���ޅ�h*᩾��1����vy��_+ �iW�	$4��W	�I?��4����(#9��ڪb��b��6b�7&��r�JM�!��:S3ޱ+wg��m��Ō�1/�1�i��α5�������le���m�C��keLc�	=H�R���	|��Q'���f���1*4�
�*�"��(oe���;��k���	��"�5�3�AVr�O{fw�5r)�됅�z�0ԙȨmi[>� (���B�5o�nyԟӁϸ�B�HJ}��ѕ���#�5�����#�-��į���e��̇�ylz7�q��f %ݣ7��r�r��}n_(�X"�XP���g� ��]N�8�	f�K�֢��R8��Q��]ψ�M���j� � �F��K �ѯ�M�M�9i�l�����,�:�/۩ɀ#�#��\�t��݀gT�bT���!p�J�v����=�J�D�@�7n�-�t����c������,&IS���1�;?�*�s�[�L׻�	-�aP�����4~�G�K�Kqݹ&p������p���/��T�j�`��9p9t��էc��af�h��zȑ���q�F)y&K��cAX�h=��$�8
��N9!�y9��}��:�p�-V���ƞ�x����<�o������'���%�i��A���y�z�\�Q��ͷ�)A�?����|������/+�T�q�K���Y��h�&O�6���Ǆ�6_u�����х1�E5����7I�Du.�ߥ^I�_�Y�,PKí�d��7�Y],��8�U� �^�`�p�����s�Y\T*�Z4�Ɨ2�.J�k�l\QOg�P��?�!�I�6:"��GD�Xu׻i%�d���ٶ�î�j|��7�͔7u��.�Nyv����$�������kS�ͩ��d��-���iL�~�H���O��s[�8��YW�9X ���C��+&���0��Ng��T,j.��Pw�K�L��M_mW�
`��tnٍ'�\J3kq��j������^� �G�@�>C�B���=�ȫ�Pi�{�ЀiL0:#SPAa+���4;���>#6fIl�7[諛)!��v؈��9��kٕF`̶����~!�f:|�:Px��ĤE�X�z�z�x��ǞRDI���&Ͳ�ˢ�T�������3�-��*i�ɺ�� 3��c��+~팏�*�>���ڕsƣ�βw��� 'c�[Y]��b\G⾲S�Q8J..�=]�����<��j��o��
ބ�8�_�%�W�ˉ�x��*��Ń��"e��o̜l���±���zg�M����n��NE���]��c�\x͜�:x�_�<@��8��s-z'��޶iN]�������6u�9�%�xn��}�TTkU� ���
Ԏu��ԃ�M��3W�Ⱦ`p'f!F5�
Kjb��=����7	fe�v<݌'��?Z�c�|�h֯�p��c^Ui���g�.k��?-�G3�,4�#�01 ҲAf>{��=o6�WyK`�*�P�jބ�C��2@�o��3�}�*g���M���]��R!��bl��q�9��s�`��Z�Ȉ���5�'�������a�$������6ŕ[� ��b��������EH�~{:�r��[��Yy�����O��}�iC���! �~�rS�G��MAk{F7�<y�T��>g�|d��%:��o�Fm{e2��B�hi!����Px��l�����l���-���Ua��g�@3 ΐ��s�.���n2o����Q�^S��9��3V( �&ƣ1��oI��+M#IʛM�p���E��>��� �{�c�K�
� >����G��S~Q��y��}I/v)r��4G��YQ�潫��l�	X�{� �;_��C03�*b��샲�,{�������4�;"ǲU5��$DWo����.2+�H��W�8�t��+����QS<���V�;sL;	����]�{O�<P=�<�=CY� ��i�h���3�5n*pseMd@ԃ�2�X)cݾKT@(h�O��V�$�GA6��?r�%�!�zgnpl��~��τ�'7	��@�AH>�� ~=t��o��B�h!v���&0F3��r?`:[���K�l]�@/`LG�����Y[�\�+
��<��t�B�BH�T�2�y��]��=y@z�7Mo�����m�l�����.��o���Z��q�t����2r����Z���@U���
P��	�sh��2	l�.�m�p�R�Ww��o�^z���ԟp`1��"\�~�����1�p�>������(ƃb	��#A���"b�x��l�[�'��v3���6��K��=����qX����So��/�9O��ѝq6���t�=�1��y�<MCWE����3������]�8�p�J`p�������#Q=���@���<�6@�yk�S�ʈf�o�\��Ya �/����nPu;c_kT�I�i���.�%��7P� �����n�j�Qe�`)$���
�i*�\*{L;rIY݌�3;iW��[���J�,�x��:��3 �@����mdK�.wX��{@W�t˩������B�&�����@�Cq�'r�v�����46*![�������zj$��K��\�g�Oz�F�G��o�
)�}4e�IdLݺŤ}<��Z��5�����2�{M`��K�p��.����܀eS��"������X|9zSD���3�|8��	z���/�|S�ݺ&��l���c������VB�����x�)0�,|НӸ�_�Xҧ�o�%�IU�����<���=t��`��£�ۑ2��~��4�!����3�T�.K�K��9��q3Fu��:)����>/�&IVځe��e��so��<Ȉ�����5����x�g�7g��	粇�أ�܅�Q�8���������s~��;YL�7y�Q��E>+��Sr��|@E��� ��Ҁ�+9���J[>N���A�G��w�U�g�/� ����P-��Ga>C\�B�f-�F\��I'49F���s�	�����J�p�~��&	FB�BۉH͐�TN��(/ˏWÔ��3�抈k�: n��� #>��)Eߟ�t�6�s���H������|�
�e4��;0I�:8��t=C��:c��������KL�:J߶��>e�&~�oߝ����P~��GYT�_��s�N���-�����CfR���'���jT�3�����Q������9�4� ƀ����>���=�u��FR�S� �{�Y$�>�>�i�N�y"C`�iv�9K�LK��"�K�h�E:>�V*��e�E������Ru�g�Q8~w^�П�����j_�qp3���^���ɧ@}g�WRV�F�
�*��>�B��"sj7p���l|���K���Q�%�5"n�$�m�uN߁� ����H�٤�md75�-?��u�2!�p���@���a�^�f/wiF4�V-戜��?���q�p����qS�L߳�rw�2��`'�*Ie��y~�[3�H�4����g�GQm��@�J�L(�A�bz_���	Fq�6P�ˋ"����d bQDv(�q�G���?��a=���a����	�YP ��܃o�l"�� �e�΋���n4�XS�?�\��7�t_2s�_&��`���'�T	�;ʇ�<+��(ve,p�ʦwK�b�d���V�>�)z;�y>���3��Rr=�z_�E莤�nJk8%����	J�Ʋ{�c�H��q�z��H� :^^0��F}	�s'ѾyEQN���Ms�V��-Yב��H�H_��y����uz@kI��,3�!���E}\��$�2��o�vY�����ވ2�p�x̩�7��p�����`�j�/OB#=m�|L����}���L"c��Do!E��$����%��al��S��nJ�՘�	G�P{�´i1�㰚[��b?ā�8M+�m|�$X�L*�<r�ގ��;���Ԕ�����2c�;$�6��"&�)������x��������f��շ�D���al`�6�˫� mr�0Zp���&KNRY��y*��e�@��?5^%��� eV8�mK��H����U�j� ��f%�E#���T��1���x�6ЙO< 3W������]U1�\�g�K8s%�+y澦�F��ky��+��x���	�1�IZd�-�O����:�����t��r�({�C�����	�H�^bD�I�ȧ�7����D�Ue���R4њLi՛�X�D�<Lp���?7�b�P��j�W��:Ͷ	G�͗��nW%ǚ�������r�)�ց,�xE�C���i�E�*ϗE�&�EQ�&�.�x��H!��* �>r����`��Jޮ���hT�����7ZP�v{%���-�Ʀ�d��-ޡZ�b�V��9p�f�B�H/�yɓu��?�D�՘2�F�pl�(zW�n���3���֐>����i���Ckt����b1�:QH;����T�qi�q�X�������W� VJ�zL�6�N���s�I�ƊjR5oq"��b���JJ���衍Zr�Y�	�l��B/l,�!�V� ���l��W�h�O�Ci.���A��#i"N�Q��`6QO���|�^�m�J&����A�n��Ix1Դ�8��|B��Ivk���VԿ ��I��i$�n�X�ħ��9�;�~�|õ��ح*�Ū�
Nh�m볊���%���%s�G�QOxB-L���Mͳ�55��-��_u�A���ف�0�X�A�3@����])����D*��`+��7Y�٣4Z�G�6��7�=���ѪtO�xT1��o�U\^%���Ia�5
Z����>G��J�-�lp�C�F�[��R����'|X��ĝb�%nb��yt�{�����/���K�G �g�Ȏ�G���r\M��>.�"!��Ρ���塐(`�J~v�����<\ԞTn����
Z⢠w�E�45^϶D��moU�f�.�R_�!޷��>�sG÷y�wQjeG��M0� �0e�ԙ����X���f,B�����/Z`�1j�:�-�r����Ēp�9���z��xb�G��a�"{�[��8iU��A,�ZS���O�Y��rƇ 9��5�"0A�q�����b7A�/B�1dtM���KO[�0��g�er�.�����:�Ӄ����,�������ϳ��K"�	��r�� v|X0NjMCd<��YRҭ�=R�Y�I}9)��8}N9]�����5��H'sU�
\�%���4��3(䨂{O�>U�<�,*����F�:qL�w��e� ކK�
\p]$����Ђ��!�2�umz�ώ5T�L�D,}� >&͍6�ʟz��Żk�I|�k!�(�='����q�;��'�l�Da�ou�i|0��3~�_vd���r�2 9�B?KcE�������ɵ^bM/�q����O�@��K�=c�\����Ȫ���[�[u�=���3�l����@�)�L)05S0���f �X>��m#�賽�Sd��9<5T
��7���?S�v7�#V&I�P�N���a<J�dJ�BL���8���͏P �g.��:Η�"�E�/��-r�xVބw��0����SN(���ż��c��贠�3^awD�s88�o�X�y�]d�y����D\��f�@���2ӑ�o���>y���<J5�:�~�v��' �.�e]���ں��2-�x������hs�[T�p题�yH��,k��%��!�^D'jU3�c�����k�/$���X�t_z�F�^_dOՋ��-ut�[����I~tJҫA�%�s�����lh�R�{'H��.�zA��{9�;׀-�U�5����3�8��/!z��=�X�	���K8=wM���-	���:庋ꬥ��S 'SM�n� �>����֑�����fk��������[���$j���XT�>�����w�*����Q'�����}(i 8�C�V����#�� ��+������C]��%�o��������
�S����"�J�*7�ƅ76�zS9f1r��r�'0���	��;�d�B�6����~�Xi�<�6�.��a����]���^+ِ��������K:n��J�ֆO�Kn�ZW}C��Ǉ#J�V/�#`�R���[�)��>L��ꚕ.<7Q��Α�0\�z &)�l��jK��\o��N�c�+n��:h �~|,� з�-���F;����M*Bm&(� $�Gb=��z�qU�DG��Rğ�/�n|� �*����-9tO]�1e�*X$8���~���̥[N��żs	�*;����Մ	T�Uo�a���u�3!6�h� ���/yc���c�~ߦͽ�=�\�>q�+v��D9Y�E���a���]�Yj���������E�i+Z�Ga4<��M�ӡ����5rQ�OR�����V�,�Wi�Z��F:5�m��e78�/�Ie�lTG�~�?Z�i\��������tY���'�P�����f�P��@>;��g��.�F�k�n	9�5�}O?ɺ����&�v��E�>�'R/���
�y�eY�� e��s2�YW���=���xf�=��:���'�E�����/)\���4(�ڏ��wN�=;�:v�53pE�}5�
�/��
��z�{��mؑ�`G3t�4H��/51� E����7-�ZHRK�VԱ�;�P���m{�ף2�U��tN��bX�e�#x%ރ8�����TQ�6��ǓF��!��T����d!�#[�l�~������4^0oœ���%"�Źeg����c�+:u��!��0V��C'l�o>�QS}�k��*�.���&�yo��̏(��%��W�U#2��V�����<F��܏�{tV}��ݠ����[=[X�%لG(�l�c����_�xD�X���@���������M��ݧ9{!������8�|�O_V�!MB�O���H�-�C�$>��y�n#;sڋ��F 6���5
�EG��%2�����G�^��L,� ��̎��~�����պ˙�i�3R��'�n[��Y��L��U�(
R�G+��(?S���z�š���V�v�|���ja�0�R��dnN��C�O�[�|��=Y5�xo��9�4�Ò;&�MӦ4g� e7`�QW�,0DT�yPHa�7�\$'�a�O1�񓈜��Iв�C@A��qՔ�	�!yO�i����U̚I����!2�+�W9<y��ǹeE�@�ar�~�a�2����3/g��2a%ꢫ錳����,,�sK}�:{�H�s��ĥs��
,�������"M������U+a�>6�z��ר�罛����b�s5^H�Jؿ�OS9�a¼x�LR�0�ԟ�<��1���-Cp$Lo�}\N �@��uY��S�q�	bt�h�oM�\�R�$�!G7^�|�`l@���^���r�ɚDf��ol�G��%�`� ���9�V�=MR��<�nK3�EǄY_9.:N�:'�$�W1�a�#�w%
�8,��H�Ff�o��mP���=i:�������S�P_���#]Ϟ�1�#N�IE}�]q������l�Jc�X�l��4��l�)]�~k��P�m�re~��	�h�؂�i���a��Z�R�"���t5+0�G<tZ(��G�X�S�L��/@\�yֹ=eK�LmJ���v��46Y����?��y?�8����o�&�ǽ��I�D�� h@C��vh�]�6�g�yQ�~���v�T�|b�1z��\�:����T(6��=��n��f-Y��$�U݊{d,u���wd�#�>�H�e��x��<�R+��(�S%�'|$��{fy10:�z�)��Ɔ�#� �c��"i�8���4R�����+Y���ZB�pʫV5
